`timescale 1ns / 1ps

module top_MH_FPGA
    (
        input clk,
        input rstn
    );

endmodule
