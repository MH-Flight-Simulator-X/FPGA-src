// Driver for the SPI communication bus between MCU and FPGA

`timescale 1ns / 1ps

module spi_driver #() ();

endmodule
